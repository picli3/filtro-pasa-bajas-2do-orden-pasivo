.title KiCad schematic
V1 /vi GND dc 10 ac 1 sin(0 10 1k 0 0)
L2 /vo_2 GND 0.6m
C1 GND /vo 10u
L1 /vi /vo 1.8m
C2 /vo_2 /vi 5.4u
.end
